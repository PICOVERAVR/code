module main_test();

reg clk = 0;
main m();

always #(1) begin
	clk <= ~clk;
end

initial begin
	
	
	
	
end
endmodule
