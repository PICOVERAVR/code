module main();
	initial begin
		$display("hello");
		$finish;
	end
endmodule
